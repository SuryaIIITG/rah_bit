`define TOTAL_APPS 1

<<<<<<< HEAD
`define PERIPLEX 0
`define GATI 1
`define MINER 2
=======
`define EXAMPLE 1

`define VERSION "1.2.0"
>>>>>>> f4d3745c2b4750be38fd7d4b5e27d7a03ac7ae14

`define GET_DATA_RAH(a) rd_data[a * RAH_PACKET_WIDTH +: RAH_PACKET_WIDTH]
`define SET_DATA_RAH(a) wr_data[a * RAH_PACKET_WIDTH +: RAH_PACKET_WIDTH]
